library verilog;
use verilog.vl_types.all;
entity Lab4_vlg_vec_tst is
end Lab4_vlg_vec_tst;
